class counter_cfg;
 static string testcase;
 static mailbox gen2bfm = new();
 static mailbox mon2cov = new();
 static virtual interface counter_if vif;
endclass
