`include "counter.sv"
`include "counter_ref.sv"
`include "interface.sv"
`include "rinterface.sv"
`include "counter_cfg.sv"
`include "counter_tx.sv"
`include "counter_gen.sv"
`include "counter_driver.sv"
`include "counter_mon.sv"
`include "counter_cov.sv"
`include "counter_scb.sv"
`include "counter_env.sv"
`include "counter_test.sv"
`include "top.sv"
